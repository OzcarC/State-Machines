`timescale 1ns/1ps

module mooreSM(input in);


endmodule