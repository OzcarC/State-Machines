`timescale 1ns/1ps

module counterDecoder(
    input stop,
);
